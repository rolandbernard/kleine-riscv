module decode (
);


endmodule
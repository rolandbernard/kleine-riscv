module memory (

);

endmodule
module core (
);


endmodule
module csr (
    input [11:0] csr_read_address,
    input csr_readable,
    input csr_writeable,
    
    input csr_write_enable,
    input [11:0] csr_write_address,
    input [11:0] csr_write_address,
    
);



endmodule
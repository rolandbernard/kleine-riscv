module fetch (

);

endmodule
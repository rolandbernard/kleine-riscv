module busio (

);


endmodule

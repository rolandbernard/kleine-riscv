module memio (

);


endmodule
module loadstore (

);

endmodule
module busio (

);


endmodule